.title KiCad schematic
.include "model/C2012X7R1E105K125AB_p.mod"
.include "model/C2012X7R2A104K125AE_p.mod"
.include "model/max976.fam"
XU2 /INP /RC VDD 0 /OUT max976
R4 /OUT 0 {RLOAD}
XU3 VDD 0 C2012X7R2A104K125AE_p
R2 /INP /OUT {RLOOP}
R1 /CTRL /INP {RIN}
R3 /RC /OUT {ROSC}
XU1 /RC 0 C2012X7R1E105K125AB_p
V1 /CTRL 0 {VCTRL}
V2 VDD 0 {VSUPPLY}
.end
